module N_bit_subtractor #(

    parameter N = 8; // N bits
) (
    input wire [N-1:0]a,
    input wire [N-1:0]b,
    input wire Cin,
    output wire [N-1:0]y,
    output wire Cout
);
    
endmodule